/scratch/nk/sram22_sky130_macros/sramgen_sram_32x32m2w8_replica_v1/sramgen_sram_32x32m2w8_replica_v1.lef