/scratch/nk/sram22_sky130_macros/sramgen_sram_512x32m4w8_replica_v1/sramgen_sram_512x32m4w8_replica_v1.lef