/home/ff/eecs151/ASAP7/asap7libs_24/techlef_misc/asap7_tech_4x_170803.lef