/scratch/nk/sram22_sky130_macros/sramgen_sram_64x32m4w32_replica_v1/sramgen_sram_64x32m4w32_replica_v1.lef