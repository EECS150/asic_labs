/scratch/nk/sram22_sky130_macros/sramgen_sram_1024x64m8w32_replica_v1/sramgen_sram_1024x64m8w32_replica_v1.lef