/scratch/nk/sram22_sky130_macros/sramgen_sram_4096x8m8w8_replica_v1/sramgen_sram_4096x8m8w8_replica_v1.lef