/home/ff/eecs151/ASAP7/asap7libs_24/lef/scaled/asap7sc7p5t_24_R_4x_170912.lef