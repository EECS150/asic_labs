`include "ALUop.vh"

module ALU(
    input [31:0] A,B,
    input [3:0] ALUop,
    output [31:0] Out
);

// Your code goes here

endmodule
